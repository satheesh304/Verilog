module SR_latch()
