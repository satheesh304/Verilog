module mux(a,s1,s2,out);
  input [3:0] a;
  input s1,s2;
  output out;

  always @(*) begin
    out=
    

  
