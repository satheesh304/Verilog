module Decoder_Tb();
  reg [1:0] a;
  wire [3:0] o;

  
