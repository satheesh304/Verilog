`include 2:1_MUX.v
`include 4:1_MUX.v

module MUX(a,s1,s2,s3,out);
output out;
input [7:0] a;
input s1,s2,s3;
wire oot1,out2;

  MUX_2X1 mux1() 
  

endmodule
