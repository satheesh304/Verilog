module N_MUX (A,S,out);
  
