module full_adder(input a, b, cin, output sum,carry);
wire w1,w2,w3;

xor(w1,a,b);
xor(sum,w1,cin);

assign w2 = a & b;
assign w3 = w1 & cin;
assign carry = w2 | w3;
endmodule

